module carry_save_adder_4_tb;
endmodule