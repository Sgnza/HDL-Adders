module not_gate(
    input wire a,
    output wire result
);

assign result = ~a;

endmodule